module top (
	input clk,    // Clock
	
);

endmodule